module test;

reg [63 : 0] first = 64'b0000000000000000000000000000000000000000000000000000000000000000;
reg [63 : 0] second = 64'b0000000000000000000000000000000000000000000000000000000000000000;

wire [64 : 0] add_result;
wire cout;

  initial begin
    $dumpfile("test.vcd");
    $dumpvars(0,test);

    # 100;
    first = 64'b0000000000000000000000000000000000000000000000000011000000010001;
    second = 64'b0000001000000000000000000000000000000000000000000010000001010000;

    # 300;
    first = 64'b0000000000000000000000110000000000011100000000000000000000010001;
    second = 64'b0000001000000000000010000000000000010000000000001011000001010000;
    
    # 500 $finish;
  end

  nbit_CLA_full_adder adder (first, second, 1'b0, add_result, cout);

  initial
     $monitor("At time %t, result = %h, cout = %b",
              $time, add_result, cout);
endmodule // test
